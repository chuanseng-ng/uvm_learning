`ifndef REGS_PKG__SV
`define REGS_PKG__SV

  package regs_pkg;

    // Import UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Reg Model UVCs

  endpackage

`endif

//End of regs_pkg
